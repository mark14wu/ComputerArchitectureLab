`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: USTC ESLAB（Embeded System Lab）
// Engineer: Haojun Xia & Xuan Wang
// Create Date: 2019/02/08
// Design Name: RISCV-Pipline CPU
// Module Name: WBSegReg
// Target Devices: Nexys4
// Tool Versions: Vivado 2017.4.1
// Description: Write Back Segment Register
//////////////////////////////////////////////////////////////////////////////////
module WBSegReg(
                input wire         clk,
                input wire         en,
                input wire         clear,
                //Data Memory Access
                input wire [31:0]  A,
                input wire [31:0]  WD,
                input wire [3:0]   WE,
                output wire [31:0] RD,
                output reg [1:0]   LoadedBytesSelect,
                //Data Memory Debug
                input wire [31:0]  A2,
                input wire [31:0]  WD2,
                input wire [3:0]   WE2,
                output wire [31:0] RD2,
                //input control signals
                input wire [31:0]  ResultM,
                output reg [31:0]  ResultW, 
                input wire [4:0]   RdM,
                output reg [4:0]   RdW,
                //output constrol signals
                input wire [2:0]   RegWriteM,
                output reg [2:0]   RegWriteW,
                input wire         MemToRegM,
                output reg         MemToRegW
                );

   //
   initial begin
      LoadedBytesSelect = 2'b00;
      RegWriteW         =  1'b0;
      MemToRegW         =  1'b0;
      ResultW           =     0;
      RdW               =  5'b0;
   end
   //
   always@(posedge clk)
     if(en)
       begin
          LoadedBytesSelect <= clear ? 2'b00 : A[1:0];
          RegWriteW         <= clear ?  1'b0 : RegWriteM;
          MemToRegW         <= clear ?  1'b0 : MemToRegM;
          ResultW           <= clear ?     0 : ResultM;
          RdW               <= clear ?  5'b0 : RdM;
       end

   wire [31:0] RD_raw;

   reg [3:0]   Wea;
   reg [31:0]   Din;

   always@(*)
     begin
        case(WE)
          4'b1111:
            begin
               Wea <= WE;
               Din <= WD;
            end
          4'b0011:
            begin
               Wea <= (A[1] == 1'b1) ? 4'b1100 : 4'b0011;
               Din <= (A[1] == 1'b1) ? {WD[15:0], 16'h0000} : {16'h0000, WD[15:0]};
            end
          4'b0001:
            begin
               Wea <= WE << A[1:0];
               Din <= WD << (A[1:0] * 8);
            end
          default:
            begin
               Wea <= 0;
               Din <= 0;
            end
        endcase // case (WE)
     end // always@ (*)

   DataRam DataRamInst (
                        .clk    (clk),                      //请补全
                        .wea    (Wea),                      //请补全
                        .addra  (A[31:2]),                      //请补全
                        .dina   (Din),                      //请补全
                        .douta  ( RD_raw         ),
                        .web    ( WE2            ),
                        .addrb  ( A2[31:2]       ),
                        .dinb   ( WD2            ),
                        .doutb  ( RD2            )
                        );
   // Add clear and stall support
   // if chip not enabled, output output last read result
   // else if chip clear, output 0
   // else output values from bram
   reg         stall_ff= 1'b0;
   reg         clear_ff= 1'b0;
   reg [31:0]  RD_old=32'b0;
   always @ (posedge clk)
     begin
        stall_ff<=~en;
        clear_ff<=clear;
        RD_old<=RD_raw;
     end

   assign RD = stall_ff ? RD_old : (clear_ff ? 32'b0 : RD_raw );

endmodule

//功能说明
//WBSegReg是Write Back段寄存器，
//类似于IDSegReg.V中对Bram的调用和拓展，它同时包含了一个同步读写的Bram
//（此处你可以调用我们提供的InstructionRam，它将会自动综合为block memory，你也可以替代性的调用xilinx的bram ip核）。
//同步读memory 相当于 异步读memory 的输出外接D触发器，需要时钟上升沿才能读取数据。
//此时如果再通过段寄存器缓存，那么需要两个时钟上升沿才能将数据传递到Ex段
//因此在段寄存器模块中调用该同步memory，直接将输出传递到WB段组合逻辑
//调用mem模块后输出为RD_raw，通过assign RD = stall_ff ? RD_old : (clear_ff ? 32'b0 : RD_raw );
//从而实现RD段寄存器stall和clear功能
//实验要求
//你需要补全上方代码，需补全的片段截取如下
//DataRam DataRamInst (
//    .clk    (???),                      //请补全
//    .wea    (???),                      //请补全
//    .addra  (???),                      //请补全
//    .dina   (???),                      //请补全
//    .douta  ( RD_raw         ),
//    .web    ( WE2            ),
//    .addrb  ( A2[31:2]       ),
//    .dinb   ( WD2            ),
//    .doutb  ( RD2            )
//);
//注意事项
//输入到DataRam的addra是字地址，一个字32bit
//请配合DataExt模块实现非字对齐字节load
//请通过补全代码实现非字对齐store
