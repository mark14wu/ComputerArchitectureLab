`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: USTC ESLAB
// Engineer: Xuan Wang (wgg@mail.ustc.edu.cn)
// 
// Create Date: 2019/02/08 16:29:41
// Design Name: RISCV-Pipline CPU
// Module Name: InstructionRamWrapper
// Target Devices: Nexys4
// Tool Versions: Vivado 2017.4.1
// Description: a Verilog-based ram which can be systhesis as BRAM
// 
//////////////////////////////////////////////////////////////////////////////////


module DataRam(
    input  clk,
    input  [ 3:0] wea, web,
    input  [31:2] addra, addrb,
    input  [31:0] dina , dinb,
    output reg [31:0] douta, doutb
);
initial begin douta=0; doutb=0; end

wire addra_valid = ( addra[31:14]==18'h0 );
wire addrb_valid = ( addrb[31:14]==18'h0 );
wire [11:0] addral = addra[13:2];
wire [11:0] addrbl = addrb[13:2];

reg [31:0] ram_cell [0:4095];

`define BTB

initial begin    // add simulation data here
    `ifdef BTB
        ram_cell[   0] = 32'h00000293;
        ram_cell[   1] = 32'h00000313;
        ram_cell[   2] = 32'h06500393;
        ram_cell[   3] = 32'h00530333;
        ram_cell[   4] = 32'h00128293;
        ram_cell[   5] = 32'hfe729ce3;
        ram_cell[   6] = 32'h00130313;
    `endif
    `ifdef BHT
        ram_cell[   0] = 32'h00000293;
        ram_cell[   1] = 32'h00000313;
        ram_cell[   2] = 32'h00000393;
        ram_cell[   3] = 32'h00a00e13;
        ram_cell[   4] = 32'h00138393;
        ram_cell[   5] = 32'h00530333;
        ram_cell[   6] = 32'h00128293;
        ram_cell[   7] = 32'hffc29ce3;
        ram_cell[   8] = 32'h00000293;
        ram_cell[   9] = 32'hffc396e3;
        ram_cell[  10] = 32'h00130313;
    
    `endif
end

always @ (posedge clk)
    douta <= addra_valid ? ram_cell[addral] : 0;
    
always @ (posedge clk)
    doutb <= addrb_valid ? ram_cell[addrbl] : 0;

always @ (posedge clk)
    if(wea[0] & addra_valid) 
        ram_cell[addral][ 7: 0] <= dina[ 7: 0];
        
always @ (posedge clk)
    if(wea[1] & addra_valid) 
        ram_cell[addral][15: 8] <= dina[15: 8];
        
always @ (posedge clk)
    if(wea[2] & addra_valid) 
        ram_cell[addral][23:16] <= dina[23:16];
        
always @ (posedge clk)
    if(wea[3] & addra_valid) 
        ram_cell[addral][31:24] <= dina[31:24];
        
always @ (posedge clk)
    if(web[0] & addrb_valid) 
        ram_cell[addrbl][ 7: 0] <= dinb[ 7: 0];
                
always @ (posedge clk)
    if(web[1] & addrb_valid) 
        ram_cell[addrbl][15: 8] <= dinb[15: 8];
                
always @ (posedge clk)
    if(web[2] & addrb_valid) 
        ram_cell[addrbl][23:16] <= dinb[23:16];
                
always @ (posedge clk)
    if(web[3] & addrb_valid) 
        ram_cell[addrbl][31:24] <= dinb[31:24];


endmodule
